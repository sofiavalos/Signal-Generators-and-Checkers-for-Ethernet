module PCS_generator
#(
    
    parameter DATA_WIDTH           = 64                                                                                                                                                                                                                                             , 
    parameter HDR_WIDTH            = 2                                                                                                                                                                                                                                              , 
    parameter FRAME_WIDTH          = DATA_WIDTH + HDR_WIDTH  /* Frame width                           */                                                                                                                                                                            ,                                                                                                                                                                                             
    parameter CONTROL_WIDTH        = 8                       /* Control width of 8 bits               */                                                                                                                                                                            ,
    parameter TRANSCODER_BLOCKS    = 4                       /* Number of transcoder blocks           */                                                                                                                                                                            ,
    parameter TRANSCODER_WIDTH     = 257                     /* Transcoder width                      */                                                                                                                                                                            ,
    parameter TRANSCODER_HDR_WIDTH = 4                       /* Transcoder header width               */                                                                                                                                                                            ,
    parameter PROB                 = 5                       /* Probability of inserting control byte */                                                                                                                                                                            
)
(
    output logic [TRANSCODER_WIDTH  - 1 : 0] o_scrambler_0   /* Output scrambler                     */                                                                                                                                                                             ,
    output logic [TRANSCODER_WIDTH  - 1 : 0] o_scrambler_1   /* Output scrambler                     */                                                                                                                                                                             ,
    output logic [TRANSCODER_WIDTH  - 1 : 0] o_transcoder_0  /* Output transcoder                    */                                                                                                                                                                             ,
    output logic [TRANSCODER_WIDTH  - 1 : 0] o_transcoder_1  /* Output transcoder                    */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_0     /* Output frame 0                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_1     /* Output frame 1                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_2     /* Output frame 2                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_3     /* Output frame 3                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_4     /* Output frame 4                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_5     /* Output frame 5                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_6     /* Output frame 6                         */                                                                                                                                                                             ,
    output logic [FRAME_WIDTH       - 1 : 0] o_frame_7     /* Output frame 7                         */                                                                                                                                                                             ,
    input  logic [TRANSCODER_BLOCKS - 1 : 0] i_data_sel_0  /* Data selector                          */                                                                                                                                                                             ,
    input  logic [TRANSCODER_BLOCKS - 1 : 0] i_data_sel_1  /* Data selector                          */                                                                                                                                                                             ,
    input  logic                             i_valid       /* Flag to enable frame generation        */                                                                                                                                                                             ,    
    input  logic                             i_random_0    /* Flag to enable random frame generation */                                                                                                                                                                             ,
    input  logic                             i_random_1    /* Flag to enable random frame generation */                                                                                                                                                                             ,
    input  logic                             i_rst_n       /* Reset                                  */                                                                                                                                                                             ,    
    input  logic                             clk           /* Clock                                  */                                                                                                                                                                             
    
);

localparam [HDR_WIDTH - 1 : 0]
    DATA_SYNC = 2'b10 /* Data sync    */                                                                                                                                                                                                                                            ,
    CTRL_SYNC = 2'b01 /* Control sync */                                                                                                                                                                                                                                            ;

localparam [CONTROL_WIDTH - 1 : 0]
    CTRL_IDLE  = 8'h00   /* Control idle     */                                                                                                                                                                                                                                     ,
    CTRL_LPI   = 8'h01   /* Control LPI      */                                                                                                                                                                                                                                     ,
    CTRL_ERROR = 8'h1E   /* Control error    */                                                                                                                                                                                                                                     ,
    CTRL_SEQ   = 8'h4B   /* Control sequence */                                                                                                                                                                                                                                     ;
    
localparam [DATA_WIDTH - 1 : 0]
    FIXED_PATTERN_0 = 64'hAAAAAAAAAAAAAAAA                                                                                                                                                                                                                                          ,
    FIXED_PATTERN_1 = 64'h3333333333333333                                                                                                                                                                                                                                          ,
    FIXED_PATTERN_2 = 64'hFFFFFFFFFFFFFFFF                                                                                                                                                                                                                                          ,
    FIXED_PATTERN_3 = 64'h0000000000000000                                                                                                                                                                                                                                          ;

localparam [CONTROL_WIDTH - 1 : 0]
    BLOCK_TYPE_FIELD_0 = 8'h1E   /* Block type field 0 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_1 = 8'h78   /* Block type field 1 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_2 = 8'h4B   /* Block type field 2 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_3 = 8'h87   /* Block type field 3 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_4 = 8'h99    /* Block type field 4 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_5 = 8'hAA   /* Block type field 5 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_6 = 8'hB4   /* Block type field 6 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_7 = 8'hCC   /* Block type field 7 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_8 = 8'hD2   /* Block type field 8 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_9 = 8'hE1   /* Block type field 9 */                                                                                                                                                                                                                           ,
    BLOCK_TYPE_FIELD_10 = 8'hF0  /* Block type field 10 */                                                                                                                                                                                                                          ;

// Local variables
logic [FRAME_WIDTH      - 1 : 0] frame_reg_0    /* Frame register */                                                                                                                                                                                                                ;
logic [FRAME_WIDTH      - 1 : 0] frame_reg_1    /* Frame register */                                                                                                                                                                                                                ;
logic [FRAME_WIDTH      - 1 : 0] frame_reg_2    /* Frame register */                                                                                                                                                                                                                ;
logic [FRAME_WIDTH      - 1 : 0] frame_reg_3    /* Frame register */                                                                                                                                                                                                                ;                                                       
logic [FRAME_WIDTH      - 1 : 0] frame_reg_4    /* Frame register */                                                                                                                                                                                                                ;
logic [FRAME_WIDTH      - 1 : 0] frame_reg_5    /* Frame register */                                                                                                                                                                                                                ;
logic [FRAME_WIDTH      - 1 : 0] frame_reg_6    /* Frame register */                                                                                                                                                                                                                ;
logic [FRAME_WIDTH      - 1 : 0] frame_reg_7    /* Frame register */                                                                                                                                                                                                                ;           
logic [TRANSCODER_WIDTH - 1 : 0] transcoder_reg_0 /* Transcoder register */                                                                                                                                                                                                         ;
logic [TRANSCODER_WIDTH - 1 : 0] transcoder_reg_1 /* Transcoder register */                                                                                                                                                                                                         ;
logic [TRANSCODER_WIDTH - 1 : 0] scrambled_data_reg_0 /* Scrambled data */                                                                                                                                                                                                          ; 
logic [TRANSCODER_WIDTH - 1 : 0] scrambled_data_reg_1 /* Scrambled data */                                                                                                                                                                                                          ;  
logic [TRANSCODER_WIDTH - 1 : 0] lfsr_value     /* Value of LFSR */                                                                                                                                                                                                                 ;

// Task to generate a PCS frame
task automatic generate_frame(
    output logic [FRAME_WIDTH - 1 : 0] o_frame      /* Output frame */                                                                                                                                                                                                              ,
    input  int                         i_number       /* Random number */                                                                                                                                                                                                             
)                                                                                                                                                                                                                                                                                   ;
    logic         [DATA_WIDTH    - 1 : 0] data_block       /* Block of data */                                                                                                                                                                                                      ; 
    logic         [CONTROL_WIDTH - 1 : 0] control_byte     /* Control byte */                                                                                                                                                                                                       ;  
    automatic int                         insert_control   /* Flag to insert control byte */                                                                                                                                                                                        ;             

    // Generate a random data block
    data_block = $urandom($time + i_number) % 64'hFFFFFFFFFFFFFFFF                                                                                                                                                                                                                  ;                                            

    // Decide wheter insert control byte or not
    insert_control = $urandom($time + i_number) % 100                                                                                                                                                                                                                               ;

    // Create the frame
    if (insert_control < PROB) begin
        // Choose a random control byte between 0 to 2
        case ($urandom($time + i_number) % 3)
            0: control_byte = CTRL_IDLE                                                                                                                                                                                                                                             ;
            1: control_byte = CTRL_LPI                                                                                                                                                                                                                                              ;
            2: control_byte = CTRL_ERROR                                                                                                                                                                                                                                            ;
        endcase
        // Choose a byte position to insert control byte
        case ($urandom($time + i_number) % 11)
            0: data_block = {BLOCK_TYPE_FIELD_0, 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            1: data_block = {BLOCK_TYPE_FIELD_1, data_block}                                                                                                                                                                                                                        ;  
            2: data_block = {BLOCK_TYPE_FIELD_2, data_block[DATA_WIDTH - 1 -:24], 4'h0, 28'h0000000}                                                                                                                                                                                ;
            3: data_block = {BLOCK_TYPE_FIELD_3, 7'b0000000                                                                                                                                                                                                                         ,
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            4: data_block = {BLOCK_TYPE_FIELD_4,  data_block[DATA_WIDTH - 1 -:08], 6'b000000                                                                                                                                                                                        ,
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            5: data_block = {BLOCK_TYPE_FIELD_5,  data_block[DATA_WIDTH - 1 -:16], 4'h0                                                                                                                                                                                             ,
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            6: data_block = {BLOCK_TYPE_FIELD_6,  data_block[DATA_WIDTH - 1 -:24], 4'h0                                                                                                                                                                                             ,
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            7: data_block = {BLOCK_TYPE_FIELD_7,  data_block[DATA_WIDTH - 1 -:32], 3'b000                                                                                                                                                                                           ,
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            8: data_block = {BLOCK_TYPE_FIELD_8,  data_block[DATA_WIDTH - 1 -:40], 2'b00                                                                                                                                                                                            ,
                             control_byte[CONTROL_WIDTH - 2 : 0]                                                                                                                                                                                                                    , 
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            9: data_block = {BLOCK_TYPE_FIELD_8,  data_block[DATA_WIDTH - 1 -:48], 2'b0                                                                                                                                                                                             ,
                             control_byte[CONTROL_WIDTH - 2 : 0]}                                                                                                                                                                                                                   ;
            10: data_block = {BLOCK_TYPE_FIELD_10, data_block[DATA_WIDTH - 1 -:56], 1'b0}                                                                                                                                                                                           ;  
        endcase
        // Use control sync if control byte is inserted
        o_frame = {CTRL_SYNC, data_block}                                                                                                                                                                                                                                           ; 
    end else begin
         // Use data sync if no control byte
        o_frame = {DATA_SYNC, data_block}                                                                                                                                                                                                                                           ;
    end
endtask

task automatic encode_frame(
    input  logic [FRAME_WIDTH - 1 : 0] frame_reg_0 /* Frame register 0 */                                                                                                                                                                                                            ,
    input  logic [FRAME_WIDTH - 1 : 0] frame_reg_1 /* Frame register 1 */                                                                                                                                                                                                            ,
    input  logic [FRAME_WIDTH - 1 : 0] frame_reg_2 /* Frame register 2 */                                                                                                                                                                                                            ,
    input  logic [FRAME_WIDTH - 1 : 0] frame_reg_3 /* Frame register 3 */                                                                                                                                                                                                            ,
    output logic[TRANSCODER_WIDTH - 1 : 0] o_transcoder
)                                                                                                                                                                                                                                                                                   ;                                      
    // transcoder output
    logic [TRANSCODER_WIDTH     - 1 : 0] transcoder                                                                                                                                                                                                                                 ; 
    // transcoder control header
    logic [TRANSCODER_HDR_WIDTH - 1 : 0] transcoder_control_hdr                                                                                                                                                                                                                     ;
    // transcoder header
    logic                                transcoder_hdr                                                                                                                                                                                                                             ;                                    
    
    // Check if the frame is a control frame
    if((frame_reg_0[FRAME_WIDTH - 1 -: 2] == DATA_SYNC) && (frame_reg_1[FRAME_WIDTH - 1 -: 2] == DATA_SYNC) && (frame_reg_2[FRAME_WIDTH - 1 -: 2] == DATA_SYNC) && (frame_reg_3[FRAME_WIDTH - 1 -: 2] == DATA_SYNC)) begin
        // Data frame with header as 1
        transcoder = {1'b1, frame_reg_0[DATA_WIDTH - 1 : 0], frame_reg_1[DATA_WIDTH - 1 : 0], frame_reg_2[DATA_WIDTH - 1 : 0], frame_reg_3[DATA_WIDTH - 1 : 0]}                                                                                                                     ;                                                                                                                                                                                                                   ;
    end
    else begin
        // Control frame with header as 0
        transcoder_hdr = 1'b0                                                                                                                                                                                                                                                       ;
        transcoder_control_hdr = {(frame_reg_0[FRAME_WIDTH - 1 -: 2] == DATA_SYNC), (frame_reg_1[FRAME_WIDTH - 1 -: 2] == DATA_SYNC), (frame_reg_2[FRAME_WIDTH - 1 -: 2] == DATA_SYNC), (frame_reg_3[FRAME_WIDTH - 1 -: 2] == DATA_SYNC)}                                           ;
        transcoder = (frame_reg_0[FRAME_WIDTH-1 -: 2] == CTRL_SYNC) ? {transcoder_hdr, transcoder_control_hdr, frame_reg_0[DATA_WIDTH - 1 -: 4], frame_reg_0[DATA_WIDTH - 9 : 0],frame_reg_1[DATA_WIDTH - 1 : 0], frame_reg_2[DATA_WIDTH - 1 : 0], frame_reg_3[DATA_WIDTH - 1 : 0]} :
                     (frame_reg_1[FRAME_WIDTH-1 -: 2] == CTRL_SYNC) ? {transcoder_hdr, transcoder_control_hdr, frame_reg_0[DATA_WIDTH - 1 : 0], frame_reg_1[DATA_WIDTH - 1 -: 4],frame_reg_1[DATA_WIDTH - 9 : 0], frame_reg_2[DATA_WIDTH - 1 : 0], frame_reg_3[DATA_WIDTH - 1 : 0]} :
                     (frame_reg_2[FRAME_WIDTH-1 -: 2] == CTRL_SYNC) ? {transcoder_hdr, transcoder_control_hdr, frame_reg_0[DATA_WIDTH - 1 : 0], frame_reg_1[DATA_WIDTH - 1 : 0],frame_reg_2[DATA_WIDTH - 1 -: 4], frame_reg_2[DATA_WIDTH - 9 : 0], frame_reg_3[DATA_WIDTH - 1 : 0]} :
                                                                      {transcoder_hdr, transcoder_control_hdr, frame_reg_0[DATA_WIDTH - 1 : 0], frame_reg_1[DATA_WIDTH - 1 : 0],frame_reg_2[DATA_WIDTH - 1 : 0], frame_reg_3[DATA_WIDTH - 1 -: 4], frame_reg_3[DATA_WIDTH - 9 : 0]} ;
    end  
    o_transcoder = transcoder                                                                                                                                                                                                                                                       ;                                                                                                                                                                                                                   ;
endtask


task automatic scrambler(        
    output logic [TRANSCODER_WIDTH - 1 : 0] scrambled_data /* Output data scrambled */                                                                                                                                                                                              ,
    input  logic [TRANSCODER_WIDTH - 1 : 0] transcoder_reg /* Input data */
)                                                                                                                                                                                                                                                                                   ;
    logic [FRAME_WIDTH - 1 : 0] data_scrambled /* Data scrambled */                                                                                                                                                                                                                 ;

    begin
        // Scrambler LFSR
        for (int i = 0; i < TRANSCODER_WIDTH; i++) begin
            data_scrambled[i] = transcoder_reg[i] ^ lfsr_value[FRAME_WIDTH - 1] /* XOR data with LFSR output */                                                                                                                                                                     ;         
            lfsr_value        = {lfsr_value[FRAME_WIDTH - 2 : 0], lfsr_value[FRAME_WIDTH] ^ lfsr_value[217] ^ lfsr_value[198]} /* Use polynomial 1 + x^39 + x^56 */                                                                                                                 ;         
        end
        // Last bit of LFSR
        data_scrambled[FRAME_WIDTH - 1] = lfsr_value[FRAME_WIDTH - 1]                                                                                                                                                                                                               ;
        // Output scrambled data
        scrambled_data = data_scrambled                                                                                                                                                                                                                                             ;            
    end

endtask


// Frame generation process
always_ff @(posedge clk or negedge i_rst_n) begin
    if (!i_rst_n) begin
        // Reset all frame registers
        frame_reg_0          <= 'b0                                                                                                                                                                                                                                                 ;                                                                                             
        frame_reg_1          <= 'b0                                                                                                                                                                                                                                                 ;                                                                                             
        frame_reg_2          <= 'b0                                                                                                                                                                                                                                                 ;                                                                                             
        frame_reg_3          <= 'b0                                                                                                                                                                                                                                                 ;
        frame_reg_4          <= 'b0                                                                                                                                                                                                                                                 ;
        frame_reg_5          <= 'b0                                                                                                                                                                                                                                                 ;
        frame_reg_6          <= 'b0                                                                                                                                                                                                                                                 ;
        frame_reg_7          <= 'b0                                                                                                                                                                                                                                                 ;
        transcoder_reg_0     <= 'b0                                                                                                                                                                                                                                                 ;                                                                                             
        transcoder_reg_1     <= 'b0                                                                                                                                                                                                                                                 ;                                                                                             
        scrambled_data_reg_0 <= 'b0                                                                                                                                                                                                                                                 ;
        scrambled_data_reg_1 <= 'b0                                                                                                                                                                                                                                                 ;
        lfsr_value           <= {TRANSCODER_WIDTH {1'b1}}                                                                                                                                                                                                                           ;
    end 
    else if(i_valid) begin
        if(i_random_0) begin
            // Generate frames for each output
            generate_frame(frame_reg_0, 043)                                                                                                                                                                                                                                        ;
            generate_frame(frame_reg_1, 086)                                                                                                                                                                                                                                        ;
            generate_frame(frame_reg_2, 127)                                                                                                                                                                                                                                        ;
            generate_frame(frame_reg_3, 065)                                                                                                                                                                                                                                        ;
       end
       else begin
            frame_reg_0 <= {((i_data_sel_0[0] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_0}                                                                                                                                                                                      ;
            frame_reg_1 <= {((i_data_sel_0[1] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_1}                                                                                                                                                                                      ;
            frame_reg_2 <= {((i_data_sel_0[2] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_2}                                                                                                                                                                                      ;
            frame_reg_3 <= {((i_data_sel_0[3] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_3}                                                                                                                                                                                      ;
       end
       if(i_random_1) begin
            generate_frame(frame_reg_4, 098)                                                                                                                                                                                                                                        ;
            generate_frame(frame_reg_5, 123)                                                                                                                                                                                                                                        ;
            generate_frame(frame_reg_6, 234)                                                                                                                                                                                                                                        ;
            generate_frame(frame_reg_7, 098)                                                                                                                                                                                                                                        ;
       end
       else begin
            frame_reg_4 <= {((i_data_sel_1[0] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_0}                                                                                                                                                                                      ;
            frame_reg_5 <= {((i_data_sel_1[1] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_1}                                                                                                                                                                                      ;
            frame_reg_6 <= {((i_data_sel_1[2] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_2}                                                                                                                                                                                      ;
            frame_reg_7 <= {((i_data_sel_1[3] == 1) ? DATA_SYNC : CTRL_SYNC), FIXED_PATTERN_3}                                                                                                                                                                                      ;
       end
       encode_frame(frame_reg_0, frame_reg_1, frame_reg_2, frame_reg_3, transcoder_reg_0)                                                                                                                                                                                           ;
       encode_frame(frame_reg_4, frame_reg_5, frame_reg_6, frame_reg_7, transcoder_reg_1)                                                                                                                                                                                           ;
       scrambler(scrambled_data_reg_0, transcoder_reg_0)                                                                                                                                                                                                                            ;
       scrambler(scrambled_data_reg_1, transcoder_reg_1)                                                                                                                                                                                                                            ;                 
    end
    else begin
        // Keep the last frame if no valid input
        frame_reg_0          <= frame_reg_0                                                                                                                                                                                                                                         ;      
        frame_reg_1          <= frame_reg_1                                                                                                                                                                                                                                         ;      
        frame_reg_2          <= frame_reg_2                                                                                                                                                                                                                                         ;      
        frame_reg_3          <= frame_reg_3                                                                                                                                                                                                                                         ;  
        frame_reg_4          <= frame_reg_4                                                                                                                                                                                                                                         ;
        frame_reg_5          <= frame_reg_5                                                                                                                                                                                                                                         ;
        frame_reg_6          <= frame_reg_6                                                                                                                                                                                                                                         ;
        frame_reg_7          <= frame_reg_7                                                                                                                                                                                                                                         ;
        transcoder_reg_0     <= transcoder_reg_0                                                                                                                                                                                                                                    ;    
        transcoder_reg_1     <= transcoder_reg_1                                                                                                                                                                                                                                    ;      
        scrambled_data_reg_0 <= scrambled_data_reg_0                                                                                                                                                                                                                                ;
        scrambled_data_reg_1 <= scrambled_data_reg_1                                                                                                                                                                                                                                ;
        lfsr_value           <= lfsr_value                                                                                                                                                                                                                                          ;
    end
end

assign o_frame_0      = frame_reg_0                                                                                                                                                                                                                                                 ;   
assign o_frame_1      = frame_reg_1                                                                                                                                                                                                                                                 ;   
assign o_frame_2      = frame_reg_2                                                                                                                                                                                                                                                 ;   
assign o_frame_3      = frame_reg_3                                                                                                                                                                                                                                                 ;   
assign o_frame_4      = frame_reg_4                                                                                                                                                                                                                                                 ;
assign o_frame_5      = frame_reg_5                                                                                                                                                                                                                                                 ;
assign o_frame_6      = frame_reg_6                                                                                                                                                                                                                                                 ;
assign o_frame_7      = frame_reg_7                                                                                                                                                                                                                                                 ;
assign o_transcoder_0 = transcoder_reg_0                                                                                                                                                                                                                                            ;
assign o_transcoder_1 = transcoder_reg_1                                                                                                                                                                                                                                            ; 
assign o_scrambler_0  = scrambled_data_reg_0                                                                                                                                                                                                                                        ;  
assign o_scrambler_1  = scrambled_data_reg_1                                                                                                                                                                                                                                        ;                                                          

endmodule
